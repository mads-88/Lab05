module circuit_b(
    // Declare inputs
    // Declare Y output
);

    // Enter logic equation here

endmodule
