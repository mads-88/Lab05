module circuit_a(
    // Declare inputs
    // Declare Y output
);

    // Enter logic equation here

endmodule
